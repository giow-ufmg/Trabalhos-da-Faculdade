module semaforo(input clk, input rst, input bt,
	output reg [2:0] A, output reg [2:0] B);
	//Insira seu codigo aqui
endmodule
